library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity RAM_1P_Demo is
	port(CLOCK50 : in std_logic;
		  KEY     : in std_logic_vector();
		  SW      : in std_logic_vector();
		  LEDR    : out std_logic_vector());
end RAM_1P_Demo;

architecture Shell of RAM_1P_Demo is
	
end Shell;